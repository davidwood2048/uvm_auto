`ifndef __${agent_name}_defines_sv__
    `define __${agent_name}_defines_sv__
//-----------------------------------------------------------------------------
// Note:
//
// ${agent_name} defines
//-----------------------------------------------------------------------------
//
// Default define for nv_small project
    `ifndef DMA_RD_REQ_PD_WIDTH
        `define DMA_RD_REQ_PD_WIDTH 48
    `endif


`define //__${agent_name}_defines_sv__
